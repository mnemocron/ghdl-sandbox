----------------------------------------------------------------------------------
-- Company:        
-- Engineer:       simon.burkhardt
-- 
-- Create Date:    2023
-- Design Name:    
-- Module Name:    
-- Project Name:   
-- Target Devices: 
-- Tool Versions:  GHDL 4.0.0
-- Description:    
-- 
-- Dependencies:   
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- this testbench acts as a streaming master, sending bursts of data
-- counting from 1-4, also asserting tlast on the 4th data packet

-- the testbench itself acts as a correct streaming master which keeps the data
-- until it is acknowledged by the DUT by asserting tready.

-- the data pattern can be influenced by the user in 2 ways
-- + Tx requests are generated by changing the pattern in p_stimuli_tready
--   the master will try to send data for as long as sim_valid_data = '1'
-- + Rx acknowledgements are generated by changing the pattern in p_stimuli_tready
--   the downstream slave after the DUT will signal ready-to-receive 
--   when sim_ready_data = '1'

-- simulate both with OPT_DATA_REG = True / False
entity tb_reset_sync is
  generic
  (
    DATA_WIDTH   : natural := 8;
    OPT_DATA_REG : boolean := True
  );
end tb_reset_sync;

architecture bh of tb_reset_sync is
  -- DUT component declaration
  component reset_deasert_sync is
    port (
      clk          : in  std_logic;
      i_resetn     : in  std_logic;
      o_resetn     : out std_logic
    );
  end component;
  
  constant CLK_PERIOD: TIME := 5 ns;

  signal clk        : std_logic;
  signal resetn     : std_logic;
  signal reset_stim : std_logic;
  signal reset_view : std_logic;

  signal clk_count : std_logic_vector(7 downto 0) := (others => '0');
begin

  -- generate clk signal
  p_clk_gen : process
  begin
   clk <= '1';
   wait for (CLK_PERIOD / 2);
   clk <= '0';
   wait for (CLK_PERIOD / 2);
   clk_count <= std_logic_vector(unsigned(clk_count) + 1);
  end process;

  -- generate ready signal
  p_stimuli : process
  begin
    reset_stim <= '1';
    wait for (CLK_PERIOD);
    wait until clk = '1';
    wait for (CLK_PERIOD/5);
    reset_stim <= '0';
    wait until clk = '1';
    wait for (CLK_PERIOD);
    wait for (CLK_PERIOD/5);
    reset_stim <= '1';
    wait for (CLK_PERIOD);
    wait for (CLK_PERIOD);
  end process;


-- DUT instance and connections
  dut_inst : reset_deasert_sync
  port map (
    clk => clk,
    i_resetn => reset_stim,
    o_resetn => reset_view
  );

end bh;
