----------------------------------------------------------------------------------
-- Company:        
-- Engineer:       simon.burkhardt
-- 
-- Create Date:    2023
-- Design Name:    
-- Module Name:    
-- Project Name:   
-- Target Devices: 
-- Tool Versions:  GHDL 4.0.0
-- Description:    
-- 
-- Dependencies:   
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
--use ieee.std_logic_arith.all;

-- this testbench acts as a streaming master, sending bursts of data
-- counting from 1-4, also asserting tlast on the 4th data packet

-- the testbench itself acts as a correct streaming master which keeps the data
-- until it is acknowledged by the DUT by asserting tready.

-- the data pattern can be influenced by the user in 2 ways
-- + Tx requests are generated by changing the pattern in p_stimuli_tready
--   the master will try to send data for as long as sim_valid_data = '1'
-- + Rx acknowledgements are generated by changing the pattern in p_stimuli_tready
--   the downstream slave after the DUT will signal ready-to-receive 
--   when sim_ready_data = '1'

-- simulate both with OPT_DATA_REG = True / False
entity tb_iir is
  generic
  (
    WIDTH_COEFFICIENTS : natural := 16;
    WIDTH_DATA         : natural := 16;
    OPT_REG_IN         : boolean := false;
    OPT_REG_OUT        : boolean := false
  );
end tb_iir;

architecture bh of tb_iir is
  -- DUT component declaration
  component iir_df1_dsp48 is
    generic (
      WIDTH_COEFFICIENTS : natural := 16;
      WIDTH_DATA         : natural := 16;
      OPT_REG_IN         : boolean := true;
      OPT_REG_OUT        : boolean := true
    );
    port (
      clk   : in  std_logic;
      d_in  : in  std_logic_vector((WIDTH_DATA-1) downto 0);
      d_out : out std_logic_vector((WIDTH_DATA-1) downto 0);
      c_a0  : in  std_logic_vector((WIDTH_COEFFICIENTS-1) downto 0);
      c_a1  : in  std_logic_vector((WIDTH_COEFFICIENTS-1) downto 0);
      c_a2  : in  std_logic_vector((WIDTH_COEFFICIENTS-1) downto 0);
      c_b0  : in  std_logic_vector((WIDTH_COEFFICIENTS-1) downto 0);
      c_b1  : in  std_logic_vector((WIDTH_COEFFICIENTS-1) downto 0)
    );
  end component;
  
  constant CLK_PERIOD: TIME := 5 ns;

  signal clk        : std_logic;
  signal resetn     : std_logic;

  signal sig_d_in  : std_logic_vector((WIDTH_DATA-1) downto 0);
  signal sig_d_out : std_logic_vector((WIDTH_DATA-1) downto 0);
  signal sig_c_a0  : std_logic_vector((WIDTH_COEFFICIENTS-1) downto 0);
  signal sig_c_a1  : std_logic_vector((WIDTH_COEFFICIENTS-1) downto 0);
  signal sig_c_a2  : std_logic_vector((WIDTH_COEFFICIENTS-1) downto 0);
  signal sig_c_b0  : std_logic_vector((WIDTH_COEFFICIENTS-1) downto 0);
  signal sig_c_b1  : std_logic_vector((WIDTH_COEFFICIENTS-1) downto 0);

  signal clk_count : std_logic_vector(7 downto 0) := (others => '0');
begin

  -- generate clk signal
  p_clk_gen : process
  begin
   clk <= '1';
   wait for (CLK_PERIOD / 2);
   clk <= '0';
   wait for (CLK_PERIOD / 2);
   clk_count <= std_logic_vector(signed(clk_count) + 1);
  end process;

  -- generate ready signal
  p_stimuli : process
  begin
    sig_c_a0 <= x"4000";
    sig_c_a1 <= x"4000";
    sig_c_a2 <= x"4000";
    sig_c_b0 <= x"0000";
    sig_c_b1 <= x"0000";
    sig_d_in <= (others => '0');
    wait until rising_edge(clk);
    sig_d_in <= x"4000";
    wait until rising_edge(clk);
    sig_d_in <= x"0000";


    wait;
  end process;


-- DUT instance and connections
  dut_inst : iir_df1_dsp48
    generic map (
      WIDTH_COEFFICIENTS => WIDTH_COEFFICIENTS,
      WIDTH_DATA         => WIDTH_DATA,
      OPT_REG_IN         => OPT_REG_IN,
      OPT_REG_OUT        => OPT_REG_OUT
    )
    port map (
      clk   => clk,
      d_in  => sig_d_in,
      d_out => sig_d_out,
      c_a0  => sig_c_a0,
      c_a1  => sig_c_a1,
      c_a2  => sig_c_a2,
      c_b0  => sig_c_b0,
      c_b1  => sig_c_b1
    );

end bh;
