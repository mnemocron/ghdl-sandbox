----------------------------------------------------------------------------------
-- Company:        
-- Engineer:       simon.burkhardt
-- 
-- Create Date:    2023-08-13
-- Design Name:    mem_sin_sfix16_2048_full 
-- Module Name:    
-- Project Name:   
-- Target Devices: Xilinx DSP48E2
-- Tool Versions:  GHDL 4.0.0-dev
-- Description:    
-- Dependencies:   
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mem_sin_sfix16_2048_full is
  generic (
    ADDR_WIDTH : natural := 11;
    DATA_WIDTH : natural := 16
  );
  port (
    a : in  std_logic_vector((ADDR_WIDTH-1) downto 0);
    o : out std_logic_vector((DATA_WIDTH-1) downto 0)
  );
end mem_sin_sfix16_2048_full;

architecture arch_imp of mem_sin_sfix16_2048_full is

  type vector_of_signed16 is array (natural range <>) of signed(15 downto 0);
  
 constant lut_data : vector_of_signed16(0 to 2047) := (
  to_signed( 16#0000#,16), to_signed( 16#0063#,16), to_signed( 16#00C7#,16), to_signed( 16#012A#,16), 
  to_signed( 16#018E#,16), to_signed( 16#01F1#,16), to_signed( 16#0255#,16), to_signed( 16#02B8#,16), 
  to_signed( 16#031C#,16), to_signed( 16#037F#,16), to_signed( 16#03E3#,16), to_signed( 16#0446#,16), 
  to_signed( 16#04AA#,16), to_signed( 16#050D#,16), to_signed( 16#0570#,16), to_signed( 16#05D4#,16), 
  to_signed( 16#0637#,16), to_signed( 16#069B#,16), to_signed( 16#06FE#,16), to_signed( 16#0761#,16), 
  to_signed( 16#07C5#,16), to_signed( 16#0828#,16), to_signed( 16#088B#,16), to_signed( 16#08EF#,16), 
  to_signed( 16#0952#,16), to_signed( 16#09B5#,16), to_signed( 16#0A18#,16), to_signed( 16#0A7C#,16), 
  to_signed( 16#0ADF#,16), to_signed( 16#0B42#,16), to_signed( 16#0BA5#,16), to_signed( 16#0C08#,16), 
  to_signed( 16#0C6B#,16), to_signed( 16#0CCE#,16), to_signed( 16#0D31#,16), to_signed( 16#0D94#,16), 
  to_signed( 16#0DF7#,16), to_signed( 16#0E5A#,16), to_signed( 16#0EBD#,16), to_signed( 16#0F20#,16), 
  to_signed( 16#0F83#,16), to_signed( 16#0FE5#,16), to_signed( 16#1048#,16), to_signed( 16#10AB#,16), 
  to_signed( 16#110D#,16), to_signed( 16#1170#,16), to_signed( 16#11D2#,16), to_signed( 16#1235#,16), 
  to_signed( 16#1297#,16), to_signed( 16#12FA#,16), to_signed( 16#135C#,16), to_signed( 16#13BF#,16), 
  to_signed( 16#1421#,16), to_signed( 16#1483#,16), to_signed( 16#14E5#,16), to_signed( 16#1547#,16), 
  to_signed( 16#15AA#,16), to_signed( 16#160C#,16), to_signed( 16#166E#,16), to_signed( 16#16D0#,16), 
  to_signed( 16#1731#,16), to_signed( 16#1793#,16), to_signed( 16#17F5#,16), to_signed( 16#1857#,16), 
  to_signed( 16#18B8#,16), to_signed( 16#191A#,16), to_signed( 16#197B#,16), to_signed( 16#19DD#,16), 
  to_signed( 16#1A3E#,16), to_signed( 16#1AA0#,16), to_signed( 16#1B01#,16), to_signed( 16#1B62#,16), 
  to_signed( 16#1BC3#,16), to_signed( 16#1C24#,16), to_signed( 16#1C85#,16), to_signed( 16#1CE6#,16), 
  to_signed( 16#1D47#,16), to_signed( 16#1DA8#,16), to_signed( 16#1E09#,16), to_signed( 16#1E69#,16), 
  to_signed( 16#1ECA#,16), to_signed( 16#1F2A#,16), to_signed( 16#1F8B#,16), to_signed( 16#1FEB#,16), 
  to_signed( 16#204B#,16), to_signed( 16#20AC#,16), to_signed( 16#210C#,16), to_signed( 16#216C#,16), 
  to_signed( 16#21CC#,16), to_signed( 16#222C#,16), to_signed( 16#228B#,16), to_signed( 16#22EB#,16), 
  to_signed( 16#234B#,16), to_signed( 16#23AA#,16), to_signed( 16#240A#,16), to_signed( 16#2469#,16), 
  to_signed( 16#24C8#,16), to_signed( 16#2528#,16), to_signed( 16#2587#,16), to_signed( 16#25E6#,16), 
  to_signed( 16#2645#,16), to_signed( 16#26A4#,16), to_signed( 16#2702#,16), to_signed( 16#2761#,16), 
  to_signed( 16#27BF#,16), to_signed( 16#281E#,16), to_signed( 16#287C#,16), to_signed( 16#28DB#,16), 
  to_signed( 16#2939#,16), to_signed( 16#2997#,16), to_signed( 16#29F5#,16), to_signed( 16#2A53#,16), 
  to_signed( 16#2AB0#,16), to_signed( 16#2B0E#,16), to_signed( 16#2B6C#,16), to_signed( 16#2BC9#,16), 
  to_signed( 16#2C26#,16), to_signed( 16#2C84#,16), to_signed( 16#2CE1#,16), to_signed( 16#2D3E#,16), 
  to_signed( 16#2D9B#,16), to_signed( 16#2DF7#,16), to_signed( 16#2E54#,16), to_signed( 16#2EB1#,16), 
  to_signed( 16#2F0D#,16), to_signed( 16#2F6A#,16), to_signed( 16#2FC6#,16), to_signed( 16#3022#,16), 
  to_signed( 16#307E#,16), to_signed( 16#30DA#,16), to_signed( 16#3136#,16), to_signed( 16#3191#,16), 
  to_signed( 16#31ED#,16), to_signed( 16#3248#,16), to_signed( 16#32A3#,16), to_signed( 16#32FF#,16), 
  to_signed( 16#335A#,16), to_signed( 16#33B5#,16), to_signed( 16#340F#,16), to_signed( 16#346A#,16), 
  to_signed( 16#34C5#,16), to_signed( 16#351F#,16), to_signed( 16#3579#,16), to_signed( 16#35D3#,16), 
  to_signed( 16#362E#,16), to_signed( 16#3687#,16), to_signed( 16#36E1#,16), to_signed( 16#373B#,16), 
  to_signed( 16#3794#,16), to_signed( 16#37EE#,16), to_signed( 16#3847#,16), to_signed( 16#38A0#,16), 
  to_signed( 16#38F9#,16), to_signed( 16#3952#,16), to_signed( 16#39AB#,16), to_signed( 16#3A03#,16), 
  to_signed( 16#3A5C#,16), to_signed( 16#3AB4#,16), to_signed( 16#3B0C#,16), to_signed( 16#3B64#,16), 
  to_signed( 16#3BBC#,16), to_signed( 16#3C13#,16), to_signed( 16#3C6B#,16), to_signed( 16#3CC2#,16), 
  to_signed( 16#3D1A#,16), to_signed( 16#3D71#,16), to_signed( 16#3DC8#,16), to_signed( 16#3E1F#,16), 
  to_signed( 16#3E75#,16), to_signed( 16#3ECC#,16), to_signed( 16#3F22#,16), to_signed( 16#3F78#,16), 
  to_signed( 16#3FCE#,16), to_signed( 16#4024#,16), to_signed( 16#407A#,16), to_signed( 16#40D0#,16), 
  to_signed( 16#4125#,16), to_signed( 16#417A#,16), to_signed( 16#41D0#,16), to_signed( 16#4225#,16), 
  to_signed( 16#4279#,16), to_signed( 16#42CE#,16), to_signed( 16#4322#,16), to_signed( 16#4377#,16), 
  to_signed( 16#43CB#,16), to_signed( 16#441F#,16), to_signed( 16#4473#,16), to_signed( 16#44C7#,16), 
  to_signed( 16#451A#,16), to_signed( 16#456D#,16), to_signed( 16#45C1#,16), to_signed( 16#4614#,16), 
  to_signed( 16#4666#,16), to_signed( 16#46B9#,16), to_signed( 16#470C#,16), to_signed( 16#475E#,16), 
  to_signed( 16#47B0#,16), to_signed( 16#4802#,16), to_signed( 16#4854#,16), to_signed( 16#48A5#,16), 
  to_signed( 16#48F7#,16), to_signed( 16#4948#,16), to_signed( 16#4999#,16), to_signed( 16#49EA#,16), 
  to_signed( 16#4A3B#,16), to_signed( 16#4A8C#,16), to_signed( 16#4ADC#,16), to_signed( 16#4B2C#,16), 
  to_signed( 16#4B7C#,16), to_signed( 16#4BCC#,16), to_signed( 16#4C1C#,16), to_signed( 16#4C6B#,16), 
  to_signed( 16#4CBA#,16), to_signed( 16#4D0A#,16), to_signed( 16#4D59#,16), to_signed( 16#4DA7#,16), 
  to_signed( 16#4DF6#,16), to_signed( 16#4E44#,16), to_signed( 16#4E92#,16), to_signed( 16#4EE0#,16), 
  to_signed( 16#4F2E#,16), to_signed( 16#4F7C#,16), to_signed( 16#4FC9#,16), to_signed( 16#5016#,16), 
  to_signed( 16#5063#,16), to_signed( 16#50B0#,16), to_signed( 16#50FD#,16), to_signed( 16#5149#,16), 
  to_signed( 16#5196#,16), to_signed( 16#51E2#,16), to_signed( 16#522E#,16), to_signed( 16#5279#,16), 
  to_signed( 16#52C5#,16), to_signed( 16#5310#,16), to_signed( 16#535B#,16), to_signed( 16#53A6#,16), 
  to_signed( 16#53F0#,16), to_signed( 16#543B#,16), to_signed( 16#5485#,16), to_signed( 16#54CF#,16), 
  to_signed( 16#5519#,16), to_signed( 16#5563#,16), to_signed( 16#55AC#,16), to_signed( 16#55F5#,16), 
  to_signed( 16#563E#,16), to_signed( 16#5687#,16), to_signed( 16#56D0#,16), to_signed( 16#5718#,16), 
  to_signed( 16#5760#,16), to_signed( 16#57A8#,16), to_signed( 16#57F0#,16), to_signed( 16#5838#,16), 
  to_signed( 16#587F#,16), to_signed( 16#58C6#,16), to_signed( 16#590D#,16), to_signed( 16#5954#,16), 
  to_signed( 16#599A#,16), to_signed( 16#59E1#,16), to_signed( 16#5A27#,16), to_signed( 16#5A6C#,16), 
  to_signed( 16#5AB2#,16), to_signed( 16#5AF7#,16), to_signed( 16#5B3D#,16), to_signed( 16#5B82#,16), 
  to_signed( 16#5BC6#,16), to_signed( 16#5C0B#,16), to_signed( 16#5C4F#,16), to_signed( 16#5C93#,16), 
  to_signed( 16#5CD7#,16), to_signed( 16#5D1B#,16), to_signed( 16#5D5E#,16), to_signed( 16#5DA1#,16), 
  to_signed( 16#5DE4#,16), to_signed( 16#5E27#,16), to_signed( 16#5E69#,16), to_signed( 16#5EAC#,16), 
  to_signed( 16#5EEE#,16), to_signed( 16#5F30#,16), to_signed( 16#5F71#,16), to_signed( 16#5FB2#,16), 
  to_signed( 16#5FF4#,16), to_signed( 16#6034#,16), to_signed( 16#6075#,16), to_signed( 16#60B6#,16), 
  to_signed( 16#60F6#,16), to_signed( 16#6136#,16), to_signed( 16#6175#,16), to_signed( 16#61B5#,16), 
  to_signed( 16#61F4#,16), to_signed( 16#6233#,16), to_signed( 16#6272#,16), to_signed( 16#62B1#,16), 
  to_signed( 16#62EF#,16), to_signed( 16#632D#,16), to_signed( 16#636B#,16), to_signed( 16#63A8#,16), 
  to_signed( 16#63E6#,16), to_signed( 16#6423#,16), to_signed( 16#6460#,16), to_signed( 16#649C#,16), 
  to_signed( 16#64D9#,16), to_signed( 16#6515#,16), to_signed( 16#6551#,16), to_signed( 16#658C#,16), 
  to_signed( 16#65C8#,16), to_signed( 16#6603#,16), to_signed( 16#663E#,16), to_signed( 16#6679#,16), 
  to_signed( 16#66B3#,16), to_signed( 16#66ED#,16), to_signed( 16#6727#,16), to_signed( 16#6761#,16), 
  to_signed( 16#679A#,16), to_signed( 16#67D3#,16), to_signed( 16#680C#,16), to_signed( 16#6845#,16), 
  to_signed( 16#687D#,16), to_signed( 16#68B6#,16), to_signed( 16#68EE#,16), to_signed( 16#6925#,16), 
  to_signed( 16#695D#,16), to_signed( 16#6994#,16), to_signed( 16#69CB#,16), to_signed( 16#6A01#,16), 
  to_signed( 16#6A38#,16), to_signed( 16#6A6E#,16), to_signed( 16#6AA4#,16), to_signed( 16#6AD9#,16), 
  to_signed( 16#6B0F#,16), to_signed( 16#6B44#,16), to_signed( 16#6B79#,16), to_signed( 16#6BAD#,16), 
  to_signed( 16#6BE2#,16), to_signed( 16#6C16#,16), to_signed( 16#6C4A#,16), to_signed( 16#6C7D#,16), 
  to_signed( 16#6CB0#,16), to_signed( 16#6CE4#,16), to_signed( 16#6D16#,16), to_signed( 16#6D49#,16), 
  to_signed( 16#6D7B#,16), to_signed( 16#6DAD#,16), to_signed( 16#6DDF#,16), to_signed( 16#6E10#,16), 
  to_signed( 16#6E41#,16), to_signed( 16#6E72#,16), to_signed( 16#6EA3#,16), to_signed( 16#6ED3#,16), 
  to_signed( 16#6F03#,16), to_signed( 16#6F33#,16), to_signed( 16#6F63#,16), to_signed( 16#6F92#,16), 
  to_signed( 16#6FC1#,16), to_signed( 16#6FF0#,16), to_signed( 16#701F#,16), to_signed( 16#704D#,16), 
  to_signed( 16#707B#,16), to_signed( 16#70A9#,16), to_signed( 16#70D6#,16), to_signed( 16#7103#,16), 
  to_signed( 16#7130#,16), to_signed( 16#715D#,16), to_signed( 16#7189#,16), to_signed( 16#71B5#,16), 
  to_signed( 16#71E1#,16), to_signed( 16#720C#,16), to_signed( 16#7238#,16), to_signed( 16#7263#,16), 
  to_signed( 16#728D#,16), to_signed( 16#72B8#,16), to_signed( 16#72E2#,16), to_signed( 16#730C#,16), 
  to_signed( 16#7335#,16), to_signed( 16#735F#,16), to_signed( 16#7388#,16), to_signed( 16#73B0#,16), 
  to_signed( 16#73D9#,16), to_signed( 16#7401#,16), to_signed( 16#7429#,16), to_signed( 16#7450#,16), 
  to_signed( 16#7478#,16), to_signed( 16#749F#,16), to_signed( 16#74C6#,16), to_signed( 16#74EC#,16), 
  to_signed( 16#7512#,16), to_signed( 16#7538#,16), to_signed( 16#755E#,16), to_signed( 16#7583#,16), 
  to_signed( 16#75A9#,16), to_signed( 16#75CD#,16), to_signed( 16#75F2#,16), to_signed( 16#7616#,16), 
  to_signed( 16#763A#,16), to_signed( 16#765E#,16), to_signed( 16#7681#,16), to_signed( 16#76A4#,16), 
  to_signed( 16#76C7#,16), to_signed( 16#76EA#,16), to_signed( 16#770C#,16), to_signed( 16#772E#,16), 
  to_signed( 16#774F#,16), to_signed( 16#7771#,16), to_signed( 16#7792#,16), to_signed( 16#77B3#,16), 
  to_signed( 16#77D3#,16), to_signed( 16#77F4#,16), to_signed( 16#7813#,16), to_signed( 16#7833#,16), 
  to_signed( 16#7852#,16), to_signed( 16#7872#,16), to_signed( 16#7890#,16), to_signed( 16#78AF#,16), 
  to_signed( 16#78CD#,16), to_signed( 16#78EB#,16), to_signed( 16#7909#,16), to_signed( 16#7926#,16), 
  to_signed( 16#7943#,16), to_signed( 16#7960#,16), to_signed( 16#797C#,16), to_signed( 16#7998#,16), 
  to_signed( 16#79B4#,16), to_signed( 16#79D0#,16), to_signed( 16#79EB#,16), to_signed( 16#7A06#,16), 
  to_signed( 16#7A21#,16), to_signed( 16#7A3B#,16), to_signed( 16#7A55#,16), to_signed( 16#7A6F#,16), 
  to_signed( 16#7A89#,16), to_signed( 16#7AA2#,16), to_signed( 16#7ABB#,16), to_signed( 16#7AD3#,16), 
  to_signed( 16#7AEC#,16), to_signed( 16#7B04#,16), to_signed( 16#7B1B#,16), to_signed( 16#7B33#,16), 
  to_signed( 16#7B4A#,16), to_signed( 16#7B61#,16), to_signed( 16#7B77#,16), to_signed( 16#7B8E#,16), 
  to_signed( 16#7BA4#,16), to_signed( 16#7BB9#,16), to_signed( 16#7BCF#,16), to_signed( 16#7BE4#,16), 
  to_signed( 16#7BF8#,16), to_signed( 16#7C0D#,16), to_signed( 16#7C21#,16), to_signed( 16#7C35#,16), 
  to_signed( 16#7C48#,16), to_signed( 16#7C5C#,16), to_signed( 16#7C6F#,16), to_signed( 16#7C81#,16), 
  to_signed( 16#7C94#,16), to_signed( 16#7CA6#,16), to_signed( 16#7CB8#,16), to_signed( 16#7CC9#,16), 
  to_signed( 16#7CDA#,16), to_signed( 16#7CEB#,16), to_signed( 16#7CFC#,16), to_signed( 16#7D0C#,16), 
  to_signed( 16#7D1C#,16), to_signed( 16#7D2C#,16), to_signed( 16#7D3B#,16), to_signed( 16#7D4A#,16), 
  to_signed( 16#7D59#,16), to_signed( 16#7D67#,16), to_signed( 16#7D75#,16), to_signed( 16#7D83#,16), 
  to_signed( 16#7D91#,16), to_signed( 16#7D9E#,16), to_signed( 16#7DAB#,16), to_signed( 16#7DB8#,16), 
  to_signed( 16#7DC4#,16), to_signed( 16#7DD0#,16), to_signed( 16#7DDC#,16), to_signed( 16#7DE7#,16), 
  to_signed( 16#7DF2#,16), to_signed( 16#7DFD#,16), to_signed( 16#7E07#,16), to_signed( 16#7E12#,16), 
  to_signed( 16#7E1C#,16), to_signed( 16#7E25#,16), to_signed( 16#7E2F#,16), to_signed( 16#7E38#,16), 
  to_signed( 16#7E40#,16), to_signed( 16#7E49#,16), to_signed( 16#7E51#,16), to_signed( 16#7E58#,16), 
  to_signed( 16#7E60#,16), to_signed( 16#7E67#,16), to_signed( 16#7E6E#,16), to_signed( 16#7E75#,16), 
  to_signed( 16#7E7B#,16), to_signed( 16#7E81#,16), to_signed( 16#7E86#,16), to_signed( 16#7E8C#,16), 
  to_signed( 16#7E91#,16), to_signed( 16#7E95#,16), to_signed( 16#7E9A#,16), to_signed( 16#7E9E#,16), 
  to_signed( 16#7EA2#,16), to_signed( 16#7EA5#,16), to_signed( 16#7EA9#,16), to_signed( 16#7EAB#,16), 
  to_signed( 16#7EAE#,16), to_signed( 16#7EB0#,16), to_signed( 16#7EB2#,16), to_signed( 16#7EB4#,16), 
  to_signed( 16#7EB5#,16), to_signed( 16#7EB6#,16), to_signed( 16#7EB7#,16), to_signed( 16#7EB8#,16), 
  to_signed( 16#7EB8#,16), to_signed( 16#7EB8#,16), to_signed( 16#7EB7#,16), to_signed( 16#7EB6#,16), 
  to_signed( 16#7EB5#,16), to_signed( 16#7EB4#,16), to_signed( 16#7EB2#,16), to_signed( 16#7EB0#,16), 
  to_signed( 16#7EAE#,16), to_signed( 16#7EAB#,16), to_signed( 16#7EA9#,16), to_signed( 16#7EA5#,16), 
  to_signed( 16#7EA2#,16), to_signed( 16#7E9E#,16), to_signed( 16#7E9A#,16), to_signed( 16#7E95#,16), 
  to_signed( 16#7E91#,16), to_signed( 16#7E8C#,16), to_signed( 16#7E86#,16), to_signed( 16#7E81#,16), 
  to_signed( 16#7E7B#,16), to_signed( 16#7E75#,16), to_signed( 16#7E6E#,16), to_signed( 16#7E67#,16), 
  to_signed( 16#7E60#,16), to_signed( 16#7E58#,16), to_signed( 16#7E51#,16), to_signed( 16#7E49#,16), 
  to_signed( 16#7E40#,16), to_signed( 16#7E38#,16), to_signed( 16#7E2F#,16), to_signed( 16#7E25#,16), 
  to_signed( 16#7E1C#,16), to_signed( 16#7E12#,16), to_signed( 16#7E07#,16), to_signed( 16#7DFD#,16), 
  to_signed( 16#7DF2#,16), to_signed( 16#7DE7#,16), to_signed( 16#7DDC#,16), to_signed( 16#7DD0#,16), 
  to_signed( 16#7DC4#,16), to_signed( 16#7DB8#,16), to_signed( 16#7DAB#,16), to_signed( 16#7D9E#,16), 
  to_signed( 16#7D91#,16), to_signed( 16#7D83#,16), to_signed( 16#7D75#,16), to_signed( 16#7D67#,16), 
  to_signed( 16#7D59#,16), to_signed( 16#7D4A#,16), to_signed( 16#7D3B#,16), to_signed( 16#7D2C#,16), 
  to_signed( 16#7D1C#,16), to_signed( 16#7D0C#,16), to_signed( 16#7CFC#,16), to_signed( 16#7CEB#,16), 
  to_signed( 16#7CDA#,16), to_signed( 16#7CC9#,16), to_signed( 16#7CB8#,16), to_signed( 16#7CA6#,16), 
  to_signed( 16#7C94#,16), to_signed( 16#7C81#,16), to_signed( 16#7C6F#,16), to_signed( 16#7C5C#,16), 
  to_signed( 16#7C48#,16), to_signed( 16#7C35#,16), to_signed( 16#7C21#,16), to_signed( 16#7C0D#,16), 
  to_signed( 16#7BF8#,16), to_signed( 16#7BE4#,16), to_signed( 16#7BCF#,16), to_signed( 16#7BB9#,16), 
  to_signed( 16#7BA4#,16), to_signed( 16#7B8E#,16), to_signed( 16#7B77#,16), to_signed( 16#7B61#,16), 
  to_signed( 16#7B4A#,16), to_signed( 16#7B33#,16), to_signed( 16#7B1B#,16), to_signed( 16#7B04#,16), 
  to_signed( 16#7AEC#,16), to_signed( 16#7AD3#,16), to_signed( 16#7ABB#,16), to_signed( 16#7AA2#,16), 
  to_signed( 16#7A89#,16), to_signed( 16#7A6F#,16), to_signed( 16#7A55#,16), to_signed( 16#7A3B#,16), 
  to_signed( 16#7A21#,16), to_signed( 16#7A06#,16), to_signed( 16#79EB#,16), to_signed( 16#79D0#,16), 
  to_signed( 16#79B4#,16), to_signed( 16#7998#,16), to_signed( 16#797C#,16), to_signed( 16#7960#,16), 
  to_signed( 16#7943#,16), to_signed( 16#7926#,16), to_signed( 16#7909#,16), to_signed( 16#78EB#,16), 
  to_signed( 16#78CD#,16), to_signed( 16#78AF#,16), to_signed( 16#7890#,16), to_signed( 16#7872#,16), 
  to_signed( 16#7852#,16), to_signed( 16#7833#,16), to_signed( 16#7813#,16), to_signed( 16#77F4#,16), 
  to_signed( 16#77D3#,16), to_signed( 16#77B3#,16), to_signed( 16#7792#,16), to_signed( 16#7771#,16), 
  to_signed( 16#774F#,16), to_signed( 16#772E#,16), to_signed( 16#770C#,16), to_signed( 16#76EA#,16), 
  to_signed( 16#76C7#,16), to_signed( 16#76A4#,16), to_signed( 16#7681#,16), to_signed( 16#765E#,16), 
  to_signed( 16#763A#,16), to_signed( 16#7616#,16), to_signed( 16#75F2#,16), to_signed( 16#75CD#,16), 
  to_signed( 16#75A9#,16), to_signed( 16#7583#,16), to_signed( 16#755E#,16), to_signed( 16#7538#,16), 
  to_signed( 16#7512#,16), to_signed( 16#74EC#,16), to_signed( 16#74C6#,16), to_signed( 16#749F#,16), 
  to_signed( 16#7478#,16), to_signed( 16#7450#,16), to_signed( 16#7429#,16), to_signed( 16#7401#,16), 
  to_signed( 16#73D9#,16), to_signed( 16#73B0#,16), to_signed( 16#7388#,16), to_signed( 16#735F#,16), 
  to_signed( 16#7335#,16), to_signed( 16#730C#,16), to_signed( 16#72E2#,16), to_signed( 16#72B8#,16), 
  to_signed( 16#728D#,16), to_signed( 16#7263#,16), to_signed( 16#7238#,16), to_signed( 16#720C#,16), 
  to_signed( 16#71E1#,16), to_signed( 16#71B5#,16), to_signed( 16#7189#,16), to_signed( 16#715D#,16), 
  to_signed( 16#7130#,16), to_signed( 16#7103#,16), to_signed( 16#70D6#,16), to_signed( 16#70A9#,16), 
  to_signed( 16#707B#,16), to_signed( 16#704D#,16), to_signed( 16#701F#,16), to_signed( 16#6FF0#,16), 
  to_signed( 16#6FC1#,16), to_signed( 16#6F92#,16), to_signed( 16#6F63#,16), to_signed( 16#6F33#,16), 
  to_signed( 16#6F03#,16), to_signed( 16#6ED3#,16), to_signed( 16#6EA3#,16), to_signed( 16#6E72#,16), 
  to_signed( 16#6E41#,16), to_signed( 16#6E10#,16), to_signed( 16#6DDF#,16), to_signed( 16#6DAD#,16), 
  to_signed( 16#6D7B#,16), to_signed( 16#6D49#,16), to_signed( 16#6D16#,16), to_signed( 16#6CE4#,16), 
  to_signed( 16#6CB0#,16), to_signed( 16#6C7D#,16), to_signed( 16#6C4A#,16), to_signed( 16#6C16#,16), 
  to_signed( 16#6BE2#,16), to_signed( 16#6BAD#,16), to_signed( 16#6B79#,16), to_signed( 16#6B44#,16), 
  to_signed( 16#6B0F#,16), to_signed( 16#6AD9#,16), to_signed( 16#6AA4#,16), to_signed( 16#6A6E#,16), 
  to_signed( 16#6A38#,16), to_signed( 16#6A01#,16), to_signed( 16#69CB#,16), to_signed( 16#6994#,16), 
  to_signed( 16#695D#,16), to_signed( 16#6925#,16), to_signed( 16#68EE#,16), to_signed( 16#68B6#,16), 
  to_signed( 16#687D#,16), to_signed( 16#6845#,16), to_signed( 16#680C#,16), to_signed( 16#67D3#,16), 
  to_signed( 16#679A#,16), to_signed( 16#6761#,16), to_signed( 16#6727#,16), to_signed( 16#66ED#,16), 
  to_signed( 16#66B3#,16), to_signed( 16#6679#,16), to_signed( 16#663E#,16), to_signed( 16#6603#,16), 
  to_signed( 16#65C8#,16), to_signed( 16#658C#,16), to_signed( 16#6551#,16), to_signed( 16#6515#,16), 
  to_signed( 16#64D9#,16), to_signed( 16#649C#,16), to_signed( 16#6460#,16), to_signed( 16#6423#,16), 
  to_signed( 16#63E6#,16), to_signed( 16#63A8#,16), to_signed( 16#636B#,16), to_signed( 16#632D#,16), 
  to_signed( 16#62EF#,16), to_signed( 16#62B1#,16), to_signed( 16#6272#,16), to_signed( 16#6233#,16), 
  to_signed( 16#61F4#,16), to_signed( 16#61B5#,16), to_signed( 16#6175#,16), to_signed( 16#6136#,16), 
  to_signed( 16#60F6#,16), to_signed( 16#60B6#,16), to_signed( 16#6075#,16), to_signed( 16#6034#,16), 
  to_signed( 16#5FF4#,16), to_signed( 16#5FB2#,16), to_signed( 16#5F71#,16), to_signed( 16#5F30#,16), 
  to_signed( 16#5EEE#,16), to_signed( 16#5EAC#,16), to_signed( 16#5E69#,16), to_signed( 16#5E27#,16), 
  to_signed( 16#5DE4#,16), to_signed( 16#5DA1#,16), to_signed( 16#5D5E#,16), to_signed( 16#5D1B#,16), 
  to_signed( 16#5CD7#,16), to_signed( 16#5C93#,16), to_signed( 16#5C4F#,16), to_signed( 16#5C0B#,16), 
  to_signed( 16#5BC6#,16), to_signed( 16#5B82#,16), to_signed( 16#5B3D#,16), to_signed( 16#5AF7#,16), 
  to_signed( 16#5AB2#,16), to_signed( 16#5A6C#,16), to_signed( 16#5A27#,16), to_signed( 16#59E1#,16), 
  to_signed( 16#599A#,16), to_signed( 16#5954#,16), to_signed( 16#590D#,16), to_signed( 16#58C6#,16), 
  to_signed( 16#587F#,16), to_signed( 16#5838#,16), to_signed( 16#57F0#,16), to_signed( 16#57A8#,16), 
  to_signed( 16#5760#,16), to_signed( 16#5718#,16), to_signed( 16#56D0#,16), to_signed( 16#5687#,16), 
  to_signed( 16#563E#,16), to_signed( 16#55F5#,16), to_signed( 16#55AC#,16), to_signed( 16#5563#,16), 
  to_signed( 16#5519#,16), to_signed( 16#54CF#,16), to_signed( 16#5485#,16), to_signed( 16#543B#,16), 
  to_signed( 16#53F0#,16), to_signed( 16#53A6#,16), to_signed( 16#535B#,16), to_signed( 16#5310#,16), 
  to_signed( 16#52C5#,16), to_signed( 16#5279#,16), to_signed( 16#522E#,16), to_signed( 16#51E2#,16), 
  to_signed( 16#5196#,16), to_signed( 16#5149#,16), to_signed( 16#50FD#,16), to_signed( 16#50B0#,16), 
  to_signed( 16#5063#,16), to_signed( 16#5016#,16), to_signed( 16#4FC9#,16), to_signed( 16#4F7C#,16), 
  to_signed( 16#4F2E#,16), to_signed( 16#4EE0#,16), to_signed( 16#4E92#,16), to_signed( 16#4E44#,16), 
  to_signed( 16#4DF6#,16), to_signed( 16#4DA7#,16), to_signed( 16#4D59#,16), to_signed( 16#4D0A#,16), 
  to_signed( 16#4CBA#,16), to_signed( 16#4C6B#,16), to_signed( 16#4C1C#,16), to_signed( 16#4BCC#,16), 
  to_signed( 16#4B7C#,16), to_signed( 16#4B2C#,16), to_signed( 16#4ADC#,16), to_signed( 16#4A8C#,16), 
  to_signed( 16#4A3B#,16), to_signed( 16#49EA#,16), to_signed( 16#4999#,16), to_signed( 16#4948#,16), 
  to_signed( 16#48F7#,16), to_signed( 16#48A5#,16), to_signed( 16#4854#,16), to_signed( 16#4802#,16), 
  to_signed( 16#47B0#,16), to_signed( 16#475E#,16), to_signed( 16#470C#,16), to_signed( 16#46B9#,16), 
  to_signed( 16#4666#,16), to_signed( 16#4614#,16), to_signed( 16#45C1#,16), to_signed( 16#456D#,16), 
  to_signed( 16#451A#,16), to_signed( 16#44C7#,16), to_signed( 16#4473#,16), to_signed( 16#441F#,16), 
  to_signed( 16#43CB#,16), to_signed( 16#4377#,16), to_signed( 16#4322#,16), to_signed( 16#42CE#,16), 
  to_signed( 16#4279#,16), to_signed( 16#4225#,16), to_signed( 16#41D0#,16), to_signed( 16#417A#,16), 
  to_signed( 16#4125#,16), to_signed( 16#40D0#,16), to_signed( 16#407A#,16), to_signed( 16#4024#,16), 
  to_signed( 16#3FCE#,16), to_signed( 16#3F78#,16), to_signed( 16#3F22#,16), to_signed( 16#3ECC#,16), 
  to_signed( 16#3E75#,16), to_signed( 16#3E1F#,16), to_signed( 16#3DC8#,16), to_signed( 16#3D71#,16), 
  to_signed( 16#3D1A#,16), to_signed( 16#3CC2#,16), to_signed( 16#3C6B#,16), to_signed( 16#3C13#,16), 
  to_signed( 16#3BBC#,16), to_signed( 16#3B64#,16), to_signed( 16#3B0C#,16), to_signed( 16#3AB4#,16), 
  to_signed( 16#3A5C#,16), to_signed( 16#3A03#,16), to_signed( 16#39AB#,16), to_signed( 16#3952#,16), 
  to_signed( 16#38F9#,16), to_signed( 16#38A0#,16), to_signed( 16#3847#,16), to_signed( 16#37EE#,16), 
  to_signed( 16#3794#,16), to_signed( 16#373B#,16), to_signed( 16#36E1#,16), to_signed( 16#3687#,16), 
  to_signed( 16#362E#,16), to_signed( 16#35D3#,16), to_signed( 16#3579#,16), to_signed( 16#351F#,16), 
  to_signed( 16#34C5#,16), to_signed( 16#346A#,16), to_signed( 16#340F#,16), to_signed( 16#33B5#,16), 
  to_signed( 16#335A#,16), to_signed( 16#32FF#,16), to_signed( 16#32A3#,16), to_signed( 16#3248#,16), 
  to_signed( 16#31ED#,16), to_signed( 16#3191#,16), to_signed( 16#3136#,16), to_signed( 16#30DA#,16), 
  to_signed( 16#307E#,16), to_signed( 16#3022#,16), to_signed( 16#2FC6#,16), to_signed( 16#2F6A#,16), 
  to_signed( 16#2F0D#,16), to_signed( 16#2EB1#,16), to_signed( 16#2E54#,16), to_signed( 16#2DF7#,16), 
  to_signed( 16#2D9B#,16), to_signed( 16#2D3E#,16), to_signed( 16#2CE1#,16), to_signed( 16#2C84#,16), 
  to_signed( 16#2C26#,16), to_signed( 16#2BC9#,16), to_signed( 16#2B6C#,16), to_signed( 16#2B0E#,16), 
  to_signed( 16#2AB0#,16), to_signed( 16#2A53#,16), to_signed( 16#29F5#,16), to_signed( 16#2997#,16), 
  to_signed( 16#2939#,16), to_signed( 16#28DB#,16), to_signed( 16#287C#,16), to_signed( 16#281E#,16), 
  to_signed( 16#27BF#,16), to_signed( 16#2761#,16), to_signed( 16#2702#,16), to_signed( 16#26A4#,16), 
  to_signed( 16#2645#,16), to_signed( 16#25E6#,16), to_signed( 16#2587#,16), to_signed( 16#2528#,16), 
  to_signed( 16#24C8#,16), to_signed( 16#2469#,16), to_signed( 16#240A#,16), to_signed( 16#23AA#,16), 
  to_signed( 16#234B#,16), to_signed( 16#22EB#,16), to_signed( 16#228B#,16), to_signed( 16#222C#,16), 
  to_signed( 16#21CC#,16), to_signed( 16#216C#,16), to_signed( 16#210C#,16), to_signed( 16#20AC#,16), 
  to_signed( 16#204B#,16), to_signed( 16#1FEB#,16), to_signed( 16#1F8B#,16), to_signed( 16#1F2A#,16), 
  to_signed( 16#1ECA#,16), to_signed( 16#1E69#,16), to_signed( 16#1E09#,16), to_signed( 16#1DA8#,16), 
  to_signed( 16#1D47#,16), to_signed( 16#1CE6#,16), to_signed( 16#1C85#,16), to_signed( 16#1C24#,16), 
  to_signed( 16#1BC3#,16), to_signed( 16#1B62#,16), to_signed( 16#1B01#,16), to_signed( 16#1AA0#,16), 
  to_signed( 16#1A3E#,16), to_signed( 16#19DD#,16), to_signed( 16#197B#,16), to_signed( 16#191A#,16), 
  to_signed( 16#18B8#,16), to_signed( 16#1857#,16), to_signed( 16#17F5#,16), to_signed( 16#1793#,16), 
  to_signed( 16#1731#,16), to_signed( 16#16D0#,16), to_signed( 16#166E#,16), to_signed( 16#160C#,16), 
  to_signed( 16#15AA#,16), to_signed( 16#1547#,16), to_signed( 16#14E5#,16), to_signed( 16#1483#,16), 
  to_signed( 16#1421#,16), to_signed( 16#13BF#,16), to_signed( 16#135C#,16), to_signed( 16#12FA#,16), 
  to_signed( 16#1297#,16), to_signed( 16#1235#,16), to_signed( 16#11D2#,16), to_signed( 16#1170#,16), 
  to_signed( 16#110D#,16), to_signed( 16#10AB#,16), to_signed( 16#1048#,16), to_signed( 16#0FE5#,16), 
  to_signed( 16#0F83#,16), to_signed( 16#0F20#,16), to_signed( 16#0EBD#,16), to_signed( 16#0E5A#,16), 
  to_signed( 16#0DF7#,16), to_signed( 16#0D94#,16), to_signed( 16#0D31#,16), to_signed( 16#0CCE#,16), 
  to_signed( 16#0C6B#,16), to_signed( 16#0C08#,16), to_signed( 16#0BA5#,16), to_signed( 16#0B42#,16), 
  to_signed( 16#0ADF#,16), to_signed( 16#0A7C#,16), to_signed( 16#0A18#,16), to_signed( 16#09B5#,16), 
  to_signed( 16#0952#,16), to_signed( 16#08EF#,16), to_signed( 16#088B#,16), to_signed( 16#0828#,16), 
  to_signed( 16#07C5#,16), to_signed( 16#0761#,16), to_signed( 16#06FE#,16), to_signed( 16#069B#,16), 
  to_signed( 16#0637#,16), to_signed( 16#05D4#,16), to_signed( 16#0570#,16), to_signed( 16#050D#,16), 
  to_signed( 16#04AA#,16), to_signed( 16#0446#,16), to_signed( 16#03E3#,16), to_signed( 16#037F#,16), 
  to_signed( 16#031C#,16), to_signed( 16#02B8#,16), to_signed( 16#0255#,16), to_signed( 16#01F1#,16), 
  to_signed( 16#018E#,16), to_signed( 16#012A#,16), to_signed( 16#00C7#,16), to_signed( 16#0063#,16), 
  to_signed( 16#0000#,16), to_signed(-16#0063#,16), to_signed(-16#00C7#,16), to_signed(-16#012A#,16), 
  to_signed(-16#018E#,16), to_signed(-16#01F1#,16), to_signed(-16#0255#,16), to_signed(-16#02B8#,16), 
  to_signed(-16#031C#,16), to_signed(-16#037F#,16), to_signed(-16#03E3#,16), to_signed(-16#0446#,16), 
  to_signed(-16#04AA#,16), to_signed(-16#050D#,16), to_signed(-16#0570#,16), to_signed(-16#05D4#,16), 
  to_signed(-16#0637#,16), to_signed(-16#069B#,16), to_signed(-16#06FE#,16), to_signed(-16#0761#,16), 
  to_signed(-16#07C5#,16), to_signed(-16#0828#,16), to_signed(-16#088B#,16), to_signed(-16#08EF#,16), 
  to_signed(-16#0952#,16), to_signed(-16#09B5#,16), to_signed(-16#0A18#,16), to_signed(-16#0A7C#,16), 
  to_signed(-16#0ADF#,16), to_signed(-16#0B42#,16), to_signed(-16#0BA5#,16), to_signed(-16#0C08#,16), 
  to_signed(-16#0C6B#,16), to_signed(-16#0CCE#,16), to_signed(-16#0D31#,16), to_signed(-16#0D94#,16), 
  to_signed(-16#0DF7#,16), to_signed(-16#0E5A#,16), to_signed(-16#0EBD#,16), to_signed(-16#0F20#,16), 
  to_signed(-16#0F83#,16), to_signed(-16#0FE5#,16), to_signed(-16#1048#,16), to_signed(-16#10AB#,16), 
  to_signed(-16#110D#,16), to_signed(-16#1170#,16), to_signed(-16#11D2#,16), to_signed(-16#1235#,16), 
  to_signed(-16#1297#,16), to_signed(-16#12FA#,16), to_signed(-16#135C#,16), to_signed(-16#13BF#,16), 
  to_signed(-16#1421#,16), to_signed(-16#1483#,16), to_signed(-16#14E5#,16), to_signed(-16#1547#,16), 
  to_signed(-16#15AA#,16), to_signed(-16#160C#,16), to_signed(-16#166E#,16), to_signed(-16#16D0#,16), 
  to_signed(-16#1731#,16), to_signed(-16#1793#,16), to_signed(-16#17F5#,16), to_signed(-16#1857#,16), 
  to_signed(-16#18B8#,16), to_signed(-16#191A#,16), to_signed(-16#197B#,16), to_signed(-16#19DD#,16), 
  to_signed(-16#1A3E#,16), to_signed(-16#1AA0#,16), to_signed(-16#1B01#,16), to_signed(-16#1B62#,16), 
  to_signed(-16#1BC3#,16), to_signed(-16#1C24#,16), to_signed(-16#1C85#,16), to_signed(-16#1CE6#,16), 
  to_signed(-16#1D47#,16), to_signed(-16#1DA8#,16), to_signed(-16#1E09#,16), to_signed(-16#1E69#,16), 
  to_signed(-16#1ECA#,16), to_signed(-16#1F2A#,16), to_signed(-16#1F8B#,16), to_signed(-16#1FEB#,16), 
  to_signed(-16#204B#,16), to_signed(-16#20AC#,16), to_signed(-16#210C#,16), to_signed(-16#216C#,16), 
  to_signed(-16#21CC#,16), to_signed(-16#222C#,16), to_signed(-16#228B#,16), to_signed(-16#22EB#,16), 
  to_signed(-16#234B#,16), to_signed(-16#23AA#,16), to_signed(-16#240A#,16), to_signed(-16#2469#,16), 
  to_signed(-16#24C8#,16), to_signed(-16#2528#,16), to_signed(-16#2587#,16), to_signed(-16#25E6#,16), 
  to_signed(-16#2645#,16), to_signed(-16#26A4#,16), to_signed(-16#2702#,16), to_signed(-16#2761#,16), 
  to_signed(-16#27BF#,16), to_signed(-16#281E#,16), to_signed(-16#287C#,16), to_signed(-16#28DB#,16), 
  to_signed(-16#2939#,16), to_signed(-16#2997#,16), to_signed(-16#29F5#,16), to_signed(-16#2A53#,16), 
  to_signed(-16#2AB0#,16), to_signed(-16#2B0E#,16), to_signed(-16#2B6C#,16), to_signed(-16#2BC9#,16), 
  to_signed(-16#2C26#,16), to_signed(-16#2C84#,16), to_signed(-16#2CE1#,16), to_signed(-16#2D3E#,16), 
  to_signed(-16#2D9B#,16), to_signed(-16#2DF7#,16), to_signed(-16#2E54#,16), to_signed(-16#2EB1#,16), 
  to_signed(-16#2F0D#,16), to_signed(-16#2F6A#,16), to_signed(-16#2FC6#,16), to_signed(-16#3022#,16), 
  to_signed(-16#307E#,16), to_signed(-16#30DA#,16), to_signed(-16#3136#,16), to_signed(-16#3191#,16), 
  to_signed(-16#31ED#,16), to_signed(-16#3248#,16), to_signed(-16#32A3#,16), to_signed(-16#32FF#,16), 
  to_signed(-16#335A#,16), to_signed(-16#33B5#,16), to_signed(-16#340F#,16), to_signed(-16#346A#,16), 
  to_signed(-16#34C5#,16), to_signed(-16#351F#,16), to_signed(-16#3579#,16), to_signed(-16#35D3#,16), 
  to_signed(-16#362E#,16), to_signed(-16#3687#,16), to_signed(-16#36E1#,16), to_signed(-16#373B#,16), 
  to_signed(-16#3794#,16), to_signed(-16#37EE#,16), to_signed(-16#3847#,16), to_signed(-16#38A0#,16), 
  to_signed(-16#38F9#,16), to_signed(-16#3952#,16), to_signed(-16#39AB#,16), to_signed(-16#3A03#,16), 
  to_signed(-16#3A5C#,16), to_signed(-16#3AB4#,16), to_signed(-16#3B0C#,16), to_signed(-16#3B64#,16), 
  to_signed(-16#3BBC#,16), to_signed(-16#3C13#,16), to_signed(-16#3C6B#,16), to_signed(-16#3CC2#,16), 
  to_signed(-16#3D1A#,16), to_signed(-16#3D71#,16), to_signed(-16#3DC8#,16), to_signed(-16#3E1F#,16), 
  to_signed(-16#3E75#,16), to_signed(-16#3ECC#,16), to_signed(-16#3F22#,16), to_signed(-16#3F78#,16), 
  to_signed(-16#3FCE#,16), to_signed(-16#4024#,16), to_signed(-16#407A#,16), to_signed(-16#40D0#,16), 
  to_signed(-16#4125#,16), to_signed(-16#417A#,16), to_signed(-16#41D0#,16), to_signed(-16#4225#,16), 
  to_signed(-16#4279#,16), to_signed(-16#42CE#,16), to_signed(-16#4322#,16), to_signed(-16#4377#,16), 
  to_signed(-16#43CB#,16), to_signed(-16#441F#,16), to_signed(-16#4473#,16), to_signed(-16#44C7#,16), 
  to_signed(-16#451A#,16), to_signed(-16#456D#,16), to_signed(-16#45C1#,16), to_signed(-16#4614#,16), 
  to_signed(-16#4666#,16), to_signed(-16#46B9#,16), to_signed(-16#470C#,16), to_signed(-16#475E#,16), 
  to_signed(-16#47B0#,16), to_signed(-16#4802#,16), to_signed(-16#4854#,16), to_signed(-16#48A5#,16), 
  to_signed(-16#48F7#,16), to_signed(-16#4948#,16), to_signed(-16#4999#,16), to_signed(-16#49EA#,16), 
  to_signed(-16#4A3B#,16), to_signed(-16#4A8C#,16), to_signed(-16#4ADC#,16), to_signed(-16#4B2C#,16), 
  to_signed(-16#4B7C#,16), to_signed(-16#4BCC#,16), to_signed(-16#4C1C#,16), to_signed(-16#4C6B#,16), 
  to_signed(-16#4CBA#,16), to_signed(-16#4D0A#,16), to_signed(-16#4D59#,16), to_signed(-16#4DA7#,16), 
  to_signed(-16#4DF6#,16), to_signed(-16#4E44#,16), to_signed(-16#4E92#,16), to_signed(-16#4EE0#,16), 
  to_signed(-16#4F2E#,16), to_signed(-16#4F7C#,16), to_signed(-16#4FC9#,16), to_signed(-16#5016#,16), 
  to_signed(-16#5063#,16), to_signed(-16#50B0#,16), to_signed(-16#50FD#,16), to_signed(-16#5149#,16), 
  to_signed(-16#5196#,16), to_signed(-16#51E2#,16), to_signed(-16#522E#,16), to_signed(-16#5279#,16), 
  to_signed(-16#52C5#,16), to_signed(-16#5310#,16), to_signed(-16#535B#,16), to_signed(-16#53A6#,16), 
  to_signed(-16#53F0#,16), to_signed(-16#543B#,16), to_signed(-16#5485#,16), to_signed(-16#54CF#,16), 
  to_signed(-16#5519#,16), to_signed(-16#5563#,16), to_signed(-16#55AC#,16), to_signed(-16#55F5#,16), 
  to_signed(-16#563E#,16), to_signed(-16#5687#,16), to_signed(-16#56D0#,16), to_signed(-16#5718#,16), 
  to_signed(-16#5760#,16), to_signed(-16#57A8#,16), to_signed(-16#57F0#,16), to_signed(-16#5838#,16), 
  to_signed(-16#587F#,16), to_signed(-16#58C6#,16), to_signed(-16#590D#,16), to_signed(-16#5954#,16), 
  to_signed(-16#599A#,16), to_signed(-16#59E1#,16), to_signed(-16#5A27#,16), to_signed(-16#5A6C#,16), 
  to_signed(-16#5AB2#,16), to_signed(-16#5AF7#,16), to_signed(-16#5B3D#,16), to_signed(-16#5B82#,16), 
  to_signed(-16#5BC6#,16), to_signed(-16#5C0B#,16), to_signed(-16#5C4F#,16), to_signed(-16#5C93#,16), 
  to_signed(-16#5CD7#,16), to_signed(-16#5D1B#,16), to_signed(-16#5D5E#,16), to_signed(-16#5DA1#,16), 
  to_signed(-16#5DE4#,16), to_signed(-16#5E27#,16), to_signed(-16#5E69#,16), to_signed(-16#5EAC#,16), 
  to_signed(-16#5EEE#,16), to_signed(-16#5F30#,16), to_signed(-16#5F71#,16), to_signed(-16#5FB2#,16), 
  to_signed(-16#5FF4#,16), to_signed(-16#6034#,16), to_signed(-16#6075#,16), to_signed(-16#60B6#,16), 
  to_signed(-16#60F6#,16), to_signed(-16#6136#,16), to_signed(-16#6175#,16), to_signed(-16#61B5#,16), 
  to_signed(-16#61F4#,16), to_signed(-16#6233#,16), to_signed(-16#6272#,16), to_signed(-16#62B1#,16), 
  to_signed(-16#62EF#,16), to_signed(-16#632D#,16), to_signed(-16#636B#,16), to_signed(-16#63A8#,16), 
  to_signed(-16#63E6#,16), to_signed(-16#6423#,16), to_signed(-16#6460#,16), to_signed(-16#649C#,16), 
  to_signed(-16#64D9#,16), to_signed(-16#6515#,16), to_signed(-16#6551#,16), to_signed(-16#658C#,16), 
  to_signed(-16#65C8#,16), to_signed(-16#6603#,16), to_signed(-16#663E#,16), to_signed(-16#6679#,16), 
  to_signed(-16#66B3#,16), to_signed(-16#66ED#,16), to_signed(-16#6727#,16), to_signed(-16#6761#,16), 
  to_signed(-16#679A#,16), to_signed(-16#67D3#,16), to_signed(-16#680C#,16), to_signed(-16#6845#,16), 
  to_signed(-16#687D#,16), to_signed(-16#68B6#,16), to_signed(-16#68EE#,16), to_signed(-16#6925#,16), 
  to_signed(-16#695D#,16), to_signed(-16#6994#,16), to_signed(-16#69CB#,16), to_signed(-16#6A01#,16), 
  to_signed(-16#6A38#,16), to_signed(-16#6A6E#,16), to_signed(-16#6AA4#,16), to_signed(-16#6AD9#,16), 
  to_signed(-16#6B0F#,16), to_signed(-16#6B44#,16), to_signed(-16#6B79#,16), to_signed(-16#6BAD#,16), 
  to_signed(-16#6BE2#,16), to_signed(-16#6C16#,16), to_signed(-16#6C4A#,16), to_signed(-16#6C7D#,16), 
  to_signed(-16#6CB0#,16), to_signed(-16#6CE4#,16), to_signed(-16#6D16#,16), to_signed(-16#6D49#,16), 
  to_signed(-16#6D7B#,16), to_signed(-16#6DAD#,16), to_signed(-16#6DDF#,16), to_signed(-16#6E10#,16), 
  to_signed(-16#6E41#,16), to_signed(-16#6E72#,16), to_signed(-16#6EA3#,16), to_signed(-16#6ED3#,16), 
  to_signed(-16#6F03#,16), to_signed(-16#6F33#,16), to_signed(-16#6F63#,16), to_signed(-16#6F92#,16), 
  to_signed(-16#6FC1#,16), to_signed(-16#6FF0#,16), to_signed(-16#701F#,16), to_signed(-16#704D#,16), 
  to_signed(-16#707B#,16), to_signed(-16#70A9#,16), to_signed(-16#70D6#,16), to_signed(-16#7103#,16), 
  to_signed(-16#7130#,16), to_signed(-16#715D#,16), to_signed(-16#7189#,16), to_signed(-16#71B5#,16), 
  to_signed(-16#71E1#,16), to_signed(-16#720C#,16), to_signed(-16#7238#,16), to_signed(-16#7263#,16), 
  to_signed(-16#728D#,16), to_signed(-16#72B8#,16), to_signed(-16#72E2#,16), to_signed(-16#730C#,16), 
  to_signed(-16#7335#,16), to_signed(-16#735F#,16), to_signed(-16#7388#,16), to_signed(-16#73B0#,16), 
  to_signed(-16#73D9#,16), to_signed(-16#7401#,16), to_signed(-16#7429#,16), to_signed(-16#7450#,16), 
  to_signed(-16#7478#,16), to_signed(-16#749F#,16), to_signed(-16#74C6#,16), to_signed(-16#74EC#,16), 
  to_signed(-16#7512#,16), to_signed(-16#7538#,16), to_signed(-16#755E#,16), to_signed(-16#7583#,16), 
  to_signed(-16#75A9#,16), to_signed(-16#75CD#,16), to_signed(-16#75F2#,16), to_signed(-16#7616#,16), 
  to_signed(-16#763A#,16), to_signed(-16#765E#,16), to_signed(-16#7681#,16), to_signed(-16#76A4#,16), 
  to_signed(-16#76C7#,16), to_signed(-16#76EA#,16), to_signed(-16#770C#,16), to_signed(-16#772E#,16), 
  to_signed(-16#774F#,16), to_signed(-16#7771#,16), to_signed(-16#7792#,16), to_signed(-16#77B3#,16), 
  to_signed(-16#77D3#,16), to_signed(-16#77F4#,16), to_signed(-16#7813#,16), to_signed(-16#7833#,16), 
  to_signed(-16#7852#,16), to_signed(-16#7872#,16), to_signed(-16#7890#,16), to_signed(-16#78AF#,16), 
  to_signed(-16#78CD#,16), to_signed(-16#78EB#,16), to_signed(-16#7909#,16), to_signed(-16#7926#,16), 
  to_signed(-16#7943#,16), to_signed(-16#7960#,16), to_signed(-16#797C#,16), to_signed(-16#7998#,16), 
  to_signed(-16#79B4#,16), to_signed(-16#79D0#,16), to_signed(-16#79EB#,16), to_signed(-16#7A06#,16), 
  to_signed(-16#7A21#,16), to_signed(-16#7A3B#,16), to_signed(-16#7A55#,16), to_signed(-16#7A6F#,16), 
  to_signed(-16#7A89#,16), to_signed(-16#7AA2#,16), to_signed(-16#7ABB#,16), to_signed(-16#7AD3#,16), 
  to_signed(-16#7AEC#,16), to_signed(-16#7B04#,16), to_signed(-16#7B1B#,16), to_signed(-16#7B33#,16), 
  to_signed(-16#7B4A#,16), to_signed(-16#7B61#,16), to_signed(-16#7B77#,16), to_signed(-16#7B8E#,16), 
  to_signed(-16#7BA4#,16), to_signed(-16#7BB9#,16), to_signed(-16#7BCF#,16), to_signed(-16#7BE4#,16), 
  to_signed(-16#7BF8#,16), to_signed(-16#7C0D#,16), to_signed(-16#7C21#,16), to_signed(-16#7C35#,16), 
  to_signed(-16#7C48#,16), to_signed(-16#7C5C#,16), to_signed(-16#7C6F#,16), to_signed(-16#7C81#,16), 
  to_signed(-16#7C94#,16), to_signed(-16#7CA6#,16), to_signed(-16#7CB8#,16), to_signed(-16#7CC9#,16), 
  to_signed(-16#7CDA#,16), to_signed(-16#7CEB#,16), to_signed(-16#7CFC#,16), to_signed(-16#7D0C#,16), 
  to_signed(-16#7D1C#,16), to_signed(-16#7D2C#,16), to_signed(-16#7D3B#,16), to_signed(-16#7D4A#,16), 
  to_signed(-16#7D59#,16), to_signed(-16#7D67#,16), to_signed(-16#7D75#,16), to_signed(-16#7D83#,16), 
  to_signed(-16#7D91#,16), to_signed(-16#7D9E#,16), to_signed(-16#7DAB#,16), to_signed(-16#7DB8#,16), 
  to_signed(-16#7DC4#,16), to_signed(-16#7DD0#,16), to_signed(-16#7DDC#,16), to_signed(-16#7DE7#,16), 
  to_signed(-16#7DF2#,16), to_signed(-16#7DFD#,16), to_signed(-16#7E07#,16), to_signed(-16#7E12#,16), 
  to_signed(-16#7E1C#,16), to_signed(-16#7E25#,16), to_signed(-16#7E2F#,16), to_signed(-16#7E38#,16), 
  to_signed(-16#7E40#,16), to_signed(-16#7E49#,16), to_signed(-16#7E51#,16), to_signed(-16#7E58#,16), 
  to_signed(-16#7E60#,16), to_signed(-16#7E67#,16), to_signed(-16#7E6E#,16), to_signed(-16#7E75#,16), 
  to_signed(-16#7E7B#,16), to_signed(-16#7E81#,16), to_signed(-16#7E86#,16), to_signed(-16#7E8C#,16), 
  to_signed(-16#7E91#,16), to_signed(-16#7E95#,16), to_signed(-16#7E9A#,16), to_signed(-16#7E9E#,16), 
  to_signed(-16#7EA2#,16), to_signed(-16#7EA5#,16), to_signed(-16#7EA9#,16), to_signed(-16#7EAB#,16), 
  to_signed(-16#7EAE#,16), to_signed(-16#7EB0#,16), to_signed(-16#7EB2#,16), to_signed(-16#7EB4#,16), 
  to_signed(-16#7EB5#,16), to_signed(-16#7EB6#,16), to_signed(-16#7EB7#,16), to_signed(-16#7EB8#,16), 
  to_signed(-16#7EB8#,16), to_signed(-16#7EB8#,16), to_signed(-16#7EB7#,16), to_signed(-16#7EB6#,16), 
  to_signed(-16#7EB5#,16), to_signed(-16#7EB4#,16), to_signed(-16#7EB2#,16), to_signed(-16#7EB0#,16), 
  to_signed(-16#7EAE#,16), to_signed(-16#7EAB#,16), to_signed(-16#7EA9#,16), to_signed(-16#7EA5#,16), 
  to_signed(-16#7EA2#,16), to_signed(-16#7E9E#,16), to_signed(-16#7E9A#,16), to_signed(-16#7E95#,16), 
  to_signed(-16#7E91#,16), to_signed(-16#7E8C#,16), to_signed(-16#7E86#,16), to_signed(-16#7E81#,16), 
  to_signed(-16#7E7B#,16), to_signed(-16#7E75#,16), to_signed(-16#7E6E#,16), to_signed(-16#7E67#,16), 
  to_signed(-16#7E60#,16), to_signed(-16#7E58#,16), to_signed(-16#7E51#,16), to_signed(-16#7E49#,16), 
  to_signed(-16#7E40#,16), to_signed(-16#7E38#,16), to_signed(-16#7E2F#,16), to_signed(-16#7E25#,16), 
  to_signed(-16#7E1C#,16), to_signed(-16#7E12#,16), to_signed(-16#7E07#,16), to_signed(-16#7DFD#,16), 
  to_signed(-16#7DF2#,16), to_signed(-16#7DE7#,16), to_signed(-16#7DDC#,16), to_signed(-16#7DD0#,16), 
  to_signed(-16#7DC4#,16), to_signed(-16#7DB8#,16), to_signed(-16#7DAB#,16), to_signed(-16#7D9E#,16), 
  to_signed(-16#7D91#,16), to_signed(-16#7D83#,16), to_signed(-16#7D75#,16), to_signed(-16#7D67#,16), 
  to_signed(-16#7D59#,16), to_signed(-16#7D4A#,16), to_signed(-16#7D3B#,16), to_signed(-16#7D2C#,16), 
  to_signed(-16#7D1C#,16), to_signed(-16#7D0C#,16), to_signed(-16#7CFC#,16), to_signed(-16#7CEB#,16), 
  to_signed(-16#7CDA#,16), to_signed(-16#7CC9#,16), to_signed(-16#7CB8#,16), to_signed(-16#7CA6#,16), 
  to_signed(-16#7C94#,16), to_signed(-16#7C81#,16), to_signed(-16#7C6F#,16), to_signed(-16#7C5C#,16), 
  to_signed(-16#7C48#,16), to_signed(-16#7C35#,16), to_signed(-16#7C21#,16), to_signed(-16#7C0D#,16), 
  to_signed(-16#7BF8#,16), to_signed(-16#7BE4#,16), to_signed(-16#7BCF#,16), to_signed(-16#7BB9#,16), 
  to_signed(-16#7BA4#,16), to_signed(-16#7B8E#,16), to_signed(-16#7B77#,16), to_signed(-16#7B61#,16), 
  to_signed(-16#7B4A#,16), to_signed(-16#7B33#,16), to_signed(-16#7B1B#,16), to_signed(-16#7B04#,16), 
  to_signed(-16#7AEC#,16), to_signed(-16#7AD3#,16), to_signed(-16#7ABB#,16), to_signed(-16#7AA2#,16), 
  to_signed(-16#7A89#,16), to_signed(-16#7A6F#,16), to_signed(-16#7A55#,16), to_signed(-16#7A3B#,16), 
  to_signed(-16#7A21#,16), to_signed(-16#7A06#,16), to_signed(-16#79EB#,16), to_signed(-16#79D0#,16), 
  to_signed(-16#79B4#,16), to_signed(-16#7998#,16), to_signed(-16#797C#,16), to_signed(-16#7960#,16), 
  to_signed(-16#7943#,16), to_signed(-16#7926#,16), to_signed(-16#7909#,16), to_signed(-16#78EB#,16), 
  to_signed(-16#78CD#,16), to_signed(-16#78AF#,16), to_signed(-16#7890#,16), to_signed(-16#7872#,16), 
  to_signed(-16#7852#,16), to_signed(-16#7833#,16), to_signed(-16#7813#,16), to_signed(-16#77F4#,16), 
  to_signed(-16#77D3#,16), to_signed(-16#77B3#,16), to_signed(-16#7792#,16), to_signed(-16#7771#,16), 
  to_signed(-16#774F#,16), to_signed(-16#772E#,16), to_signed(-16#770C#,16), to_signed(-16#76EA#,16), 
  to_signed(-16#76C7#,16), to_signed(-16#76A4#,16), to_signed(-16#7681#,16), to_signed(-16#765E#,16), 
  to_signed(-16#763A#,16), to_signed(-16#7616#,16), to_signed(-16#75F2#,16), to_signed(-16#75CD#,16), 
  to_signed(-16#75A9#,16), to_signed(-16#7583#,16), to_signed(-16#755E#,16), to_signed(-16#7538#,16), 
  to_signed(-16#7512#,16), to_signed(-16#74EC#,16), to_signed(-16#74C6#,16), to_signed(-16#749F#,16), 
  to_signed(-16#7478#,16), to_signed(-16#7450#,16), to_signed(-16#7429#,16), to_signed(-16#7401#,16), 
  to_signed(-16#73D9#,16), to_signed(-16#73B0#,16), to_signed(-16#7388#,16), to_signed(-16#735F#,16), 
  to_signed(-16#7335#,16), to_signed(-16#730C#,16), to_signed(-16#72E2#,16), to_signed(-16#72B8#,16), 
  to_signed(-16#728D#,16), to_signed(-16#7263#,16), to_signed(-16#7238#,16), to_signed(-16#720C#,16), 
  to_signed(-16#71E1#,16), to_signed(-16#71B5#,16), to_signed(-16#7189#,16), to_signed(-16#715D#,16), 
  to_signed(-16#7130#,16), to_signed(-16#7103#,16), to_signed(-16#70D6#,16), to_signed(-16#70A9#,16), 
  to_signed(-16#707B#,16), to_signed(-16#704D#,16), to_signed(-16#701F#,16), to_signed(-16#6FF0#,16), 
  to_signed(-16#6FC1#,16), to_signed(-16#6F92#,16), to_signed(-16#6F63#,16), to_signed(-16#6F33#,16), 
  to_signed(-16#6F03#,16), to_signed(-16#6ED3#,16), to_signed(-16#6EA3#,16), to_signed(-16#6E72#,16), 
  to_signed(-16#6E41#,16), to_signed(-16#6E10#,16), to_signed(-16#6DDF#,16), to_signed(-16#6DAD#,16), 
  to_signed(-16#6D7B#,16), to_signed(-16#6D49#,16), to_signed(-16#6D16#,16), to_signed(-16#6CE4#,16), 
  to_signed(-16#6CB0#,16), to_signed(-16#6C7D#,16), to_signed(-16#6C4A#,16), to_signed(-16#6C16#,16), 
  to_signed(-16#6BE2#,16), to_signed(-16#6BAD#,16), to_signed(-16#6B79#,16), to_signed(-16#6B44#,16), 
  to_signed(-16#6B0F#,16), to_signed(-16#6AD9#,16), to_signed(-16#6AA4#,16), to_signed(-16#6A6E#,16), 
  to_signed(-16#6A38#,16), to_signed(-16#6A01#,16), to_signed(-16#69CB#,16), to_signed(-16#6994#,16), 
  to_signed(-16#695D#,16), to_signed(-16#6925#,16), to_signed(-16#68EE#,16), to_signed(-16#68B6#,16), 
  to_signed(-16#687D#,16), to_signed(-16#6845#,16), to_signed(-16#680C#,16), to_signed(-16#67D3#,16), 
  to_signed(-16#679A#,16), to_signed(-16#6761#,16), to_signed(-16#6727#,16), to_signed(-16#66ED#,16), 
  to_signed(-16#66B3#,16), to_signed(-16#6679#,16), to_signed(-16#663E#,16), to_signed(-16#6603#,16), 
  to_signed(-16#65C8#,16), to_signed(-16#658C#,16), to_signed(-16#6551#,16), to_signed(-16#6515#,16), 
  to_signed(-16#64D9#,16), to_signed(-16#649C#,16), to_signed(-16#6460#,16), to_signed(-16#6423#,16), 
  to_signed(-16#63E6#,16), to_signed(-16#63A8#,16), to_signed(-16#636B#,16), to_signed(-16#632D#,16), 
  to_signed(-16#62EF#,16), to_signed(-16#62B1#,16), to_signed(-16#6272#,16), to_signed(-16#6233#,16), 
  to_signed(-16#61F4#,16), to_signed(-16#61B5#,16), to_signed(-16#6175#,16), to_signed(-16#6136#,16), 
  to_signed(-16#60F6#,16), to_signed(-16#60B6#,16), to_signed(-16#6075#,16), to_signed(-16#6034#,16), 
  to_signed(-16#5FF4#,16), to_signed(-16#5FB2#,16), to_signed(-16#5F71#,16), to_signed(-16#5F30#,16), 
  to_signed(-16#5EEE#,16), to_signed(-16#5EAC#,16), to_signed(-16#5E69#,16), to_signed(-16#5E27#,16), 
  to_signed(-16#5DE4#,16), to_signed(-16#5DA1#,16), to_signed(-16#5D5E#,16), to_signed(-16#5D1B#,16), 
  to_signed(-16#5CD7#,16), to_signed(-16#5C93#,16), to_signed(-16#5C4F#,16), to_signed(-16#5C0B#,16), 
  to_signed(-16#5BC6#,16), to_signed(-16#5B82#,16), to_signed(-16#5B3D#,16), to_signed(-16#5AF7#,16), 
  to_signed(-16#5AB2#,16), to_signed(-16#5A6C#,16), to_signed(-16#5A27#,16), to_signed(-16#59E1#,16), 
  to_signed(-16#599A#,16), to_signed(-16#5954#,16), to_signed(-16#590D#,16), to_signed(-16#58C6#,16), 
  to_signed(-16#587F#,16), to_signed(-16#5838#,16), to_signed(-16#57F0#,16), to_signed(-16#57A8#,16), 
  to_signed(-16#5760#,16), to_signed(-16#5718#,16), to_signed(-16#56D0#,16), to_signed(-16#5687#,16), 
  to_signed(-16#563E#,16), to_signed(-16#55F5#,16), to_signed(-16#55AC#,16), to_signed(-16#5563#,16), 
  to_signed(-16#5519#,16), to_signed(-16#54CF#,16), to_signed(-16#5485#,16), to_signed(-16#543B#,16), 
  to_signed(-16#53F0#,16), to_signed(-16#53A6#,16), to_signed(-16#535B#,16), to_signed(-16#5310#,16), 
  to_signed(-16#52C5#,16), to_signed(-16#5279#,16), to_signed(-16#522E#,16), to_signed(-16#51E2#,16), 
  to_signed(-16#5196#,16), to_signed(-16#5149#,16), to_signed(-16#50FD#,16), to_signed(-16#50B0#,16), 
  to_signed(-16#5063#,16), to_signed(-16#5016#,16), to_signed(-16#4FC9#,16), to_signed(-16#4F7C#,16), 
  to_signed(-16#4F2E#,16), to_signed(-16#4EE0#,16), to_signed(-16#4E92#,16), to_signed(-16#4E44#,16), 
  to_signed(-16#4DF6#,16), to_signed(-16#4DA7#,16), to_signed(-16#4D59#,16), to_signed(-16#4D0A#,16), 
  to_signed(-16#4CBA#,16), to_signed(-16#4C6B#,16), to_signed(-16#4C1C#,16), to_signed(-16#4BCC#,16), 
  to_signed(-16#4B7C#,16), to_signed(-16#4B2C#,16), to_signed(-16#4ADC#,16), to_signed(-16#4A8C#,16), 
  to_signed(-16#4A3B#,16), to_signed(-16#49EA#,16), to_signed(-16#4999#,16), to_signed(-16#4948#,16), 
  to_signed(-16#48F7#,16), to_signed(-16#48A5#,16), to_signed(-16#4854#,16), to_signed(-16#4802#,16), 
  to_signed(-16#47B0#,16), to_signed(-16#475E#,16), to_signed(-16#470C#,16), to_signed(-16#46B9#,16), 
  to_signed(-16#4666#,16), to_signed(-16#4614#,16), to_signed(-16#45C1#,16), to_signed(-16#456D#,16), 
  to_signed(-16#451A#,16), to_signed(-16#44C7#,16), to_signed(-16#4473#,16), to_signed(-16#441F#,16), 
  to_signed(-16#43CB#,16), to_signed(-16#4377#,16), to_signed(-16#4322#,16), to_signed(-16#42CE#,16), 
  to_signed(-16#4279#,16), to_signed(-16#4225#,16), to_signed(-16#41D0#,16), to_signed(-16#417A#,16), 
  to_signed(-16#4125#,16), to_signed(-16#40D0#,16), to_signed(-16#407A#,16), to_signed(-16#4024#,16), 
  to_signed(-16#3FCE#,16), to_signed(-16#3F78#,16), to_signed(-16#3F22#,16), to_signed(-16#3ECC#,16), 
  to_signed(-16#3E75#,16), to_signed(-16#3E1F#,16), to_signed(-16#3DC8#,16), to_signed(-16#3D71#,16), 
  to_signed(-16#3D1A#,16), to_signed(-16#3CC2#,16), to_signed(-16#3C6B#,16), to_signed(-16#3C13#,16), 
  to_signed(-16#3BBC#,16), to_signed(-16#3B64#,16), to_signed(-16#3B0C#,16), to_signed(-16#3AB4#,16), 
  to_signed(-16#3A5C#,16), to_signed(-16#3A03#,16), to_signed(-16#39AB#,16), to_signed(-16#3952#,16), 
  to_signed(-16#38F9#,16), to_signed(-16#38A0#,16), to_signed(-16#3847#,16), to_signed(-16#37EE#,16), 
  to_signed(-16#3794#,16), to_signed(-16#373B#,16), to_signed(-16#36E1#,16), to_signed(-16#3687#,16), 
  to_signed(-16#362E#,16), to_signed(-16#35D3#,16), to_signed(-16#3579#,16), to_signed(-16#351F#,16), 
  to_signed(-16#34C5#,16), to_signed(-16#346A#,16), to_signed(-16#340F#,16), to_signed(-16#33B5#,16), 
  to_signed(-16#335A#,16), to_signed(-16#32FF#,16), to_signed(-16#32A3#,16), to_signed(-16#3248#,16), 
  to_signed(-16#31ED#,16), to_signed(-16#3191#,16), to_signed(-16#3136#,16), to_signed(-16#30DA#,16), 
  to_signed(-16#307E#,16), to_signed(-16#3022#,16), to_signed(-16#2FC6#,16), to_signed(-16#2F6A#,16), 
  to_signed(-16#2F0D#,16), to_signed(-16#2EB1#,16), to_signed(-16#2E54#,16), to_signed(-16#2DF7#,16), 
  to_signed(-16#2D9B#,16), to_signed(-16#2D3E#,16), to_signed(-16#2CE1#,16), to_signed(-16#2C84#,16), 
  to_signed(-16#2C26#,16), to_signed(-16#2BC9#,16), to_signed(-16#2B6C#,16), to_signed(-16#2B0E#,16), 
  to_signed(-16#2AB0#,16), to_signed(-16#2A53#,16), to_signed(-16#29F5#,16), to_signed(-16#2997#,16), 
  to_signed(-16#2939#,16), to_signed(-16#28DB#,16), to_signed(-16#287C#,16), to_signed(-16#281E#,16), 
  to_signed(-16#27BF#,16), to_signed(-16#2761#,16), to_signed(-16#2702#,16), to_signed(-16#26A4#,16), 
  to_signed(-16#2645#,16), to_signed(-16#25E6#,16), to_signed(-16#2587#,16), to_signed(-16#2528#,16), 
  to_signed(-16#24C8#,16), to_signed(-16#2469#,16), to_signed(-16#240A#,16), to_signed(-16#23AA#,16), 
  to_signed(-16#234B#,16), to_signed(-16#22EB#,16), to_signed(-16#228B#,16), to_signed(-16#222C#,16), 
  to_signed(-16#21CC#,16), to_signed(-16#216C#,16), to_signed(-16#210C#,16), to_signed(-16#20AC#,16), 
  to_signed(-16#204B#,16), to_signed(-16#1FEB#,16), to_signed(-16#1F8B#,16), to_signed(-16#1F2A#,16), 
  to_signed(-16#1ECA#,16), to_signed(-16#1E69#,16), to_signed(-16#1E09#,16), to_signed(-16#1DA8#,16), 
  to_signed(-16#1D47#,16), to_signed(-16#1CE6#,16), to_signed(-16#1C85#,16), to_signed(-16#1C24#,16), 
  to_signed(-16#1BC3#,16), to_signed(-16#1B62#,16), to_signed(-16#1B01#,16), to_signed(-16#1AA0#,16), 
  to_signed(-16#1A3E#,16), to_signed(-16#19DD#,16), to_signed(-16#197B#,16), to_signed(-16#191A#,16), 
  to_signed(-16#18B8#,16), to_signed(-16#1857#,16), to_signed(-16#17F5#,16), to_signed(-16#1793#,16), 
  to_signed(-16#1731#,16), to_signed(-16#16D0#,16), to_signed(-16#166E#,16), to_signed(-16#160C#,16), 
  to_signed(-16#15AA#,16), to_signed(-16#1547#,16), to_signed(-16#14E5#,16), to_signed(-16#1483#,16), 
  to_signed(-16#1421#,16), to_signed(-16#13BF#,16), to_signed(-16#135C#,16), to_signed(-16#12FA#,16), 
  to_signed(-16#1297#,16), to_signed(-16#1235#,16), to_signed(-16#11D2#,16), to_signed(-16#1170#,16), 
  to_signed(-16#110D#,16), to_signed(-16#10AB#,16), to_signed(-16#1048#,16), to_signed(-16#0FE5#,16), 
  to_signed(-16#0F83#,16), to_signed(-16#0F20#,16), to_signed(-16#0EBD#,16), to_signed(-16#0E5A#,16), 
  to_signed(-16#0DF7#,16), to_signed(-16#0D94#,16), to_signed(-16#0D31#,16), to_signed(-16#0CCE#,16), 
  to_signed(-16#0C6B#,16), to_signed(-16#0C08#,16), to_signed(-16#0BA5#,16), to_signed(-16#0B42#,16), 
  to_signed(-16#0ADF#,16), to_signed(-16#0A7C#,16), to_signed(-16#0A18#,16), to_signed(-16#09B5#,16), 
  to_signed(-16#0952#,16), to_signed(-16#08EF#,16), to_signed(-16#088B#,16), to_signed(-16#0828#,16), 
  to_signed(-16#07C5#,16), to_signed(-16#0761#,16), to_signed(-16#06FE#,16), to_signed(-16#069B#,16), 
  to_signed(-16#0637#,16), to_signed(-16#05D4#,16), to_signed(-16#0570#,16), to_signed(-16#050D#,16), 
  to_signed(-16#04AA#,16), to_signed(-16#0446#,16), to_signed(-16#03E3#,16), to_signed(-16#037F#,16), 
  to_signed(-16#031C#,16), to_signed(-16#02B8#,16), to_signed(-16#0255#,16), to_signed(-16#01F1#,16), 
  to_signed(-16#018E#,16), to_signed(-16#012A#,16), to_signed(-16#00C7#,16), to_signed(-16#0063#,16)
);

  signal selector : unsigned((ADDR_WIDTH-1) downto 0) := (others => '0');
begin
  selector <= unsigned(a);
  o <= std_logic_vector(lut_data(to_integer(selector)));

end arch_imp;
